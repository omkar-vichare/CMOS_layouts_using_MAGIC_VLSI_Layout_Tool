magic
tech sky130A
timestamp 1734980426
<< nwell >>
rect -545 -20 610 240
<< nmos >>
rect -475 -295 -460 -240
rect -410 -295 -395 -240
rect -180 -295 -165 -185
rect 25 -295 40 -185
rect 90 -295 105 -185
rect 235 -295 250 -185
rect 300 -295 315 -185
rect 485 -295 500 -185
<< pmos >>
rect -475 0 -460 220
rect -410 0 -395 220
rect -160 0 -145 220
rect 25 0 40 220
rect 90 0 105 220
rect 235 0 250 220
rect 300 0 315 220
rect 485 0 500 220
<< ndiff >>
rect -225 -195 -180 -185
rect -225 -230 -215 -195
rect -195 -230 -180 -195
rect -525 -250 -475 -240
rect -525 -285 -510 -250
rect -490 -285 -475 -250
rect -525 -295 -475 -285
rect -460 -250 -410 -240
rect -460 -285 -445 -250
rect -425 -285 -410 -250
rect -460 -295 -410 -285
rect -395 -250 -350 -240
rect -395 -285 -380 -250
rect -360 -285 -350 -250
rect -395 -295 -350 -285
rect -225 -250 -180 -230
rect -225 -285 -215 -250
rect -195 -285 -180 -250
rect -225 -295 -180 -285
rect -165 -195 -115 -185
rect -165 -230 -150 -195
rect -130 -230 -115 -195
rect -165 -250 -115 -230
rect -165 -285 -150 -250
rect -130 -285 -115 -250
rect -165 -295 -115 -285
rect -25 -195 25 -185
rect -25 -230 -10 -195
rect 10 -230 25 -195
rect -25 -250 25 -230
rect -25 -285 -10 -250
rect 10 -285 25 -250
rect -25 -295 25 -285
rect 40 -195 90 -185
rect 40 -230 55 -195
rect 75 -230 90 -195
rect 40 -250 90 -230
rect 40 -285 55 -250
rect 75 -285 90 -250
rect 40 -295 90 -285
rect 105 -195 155 -185
rect 105 -230 120 -195
rect 140 -230 155 -195
rect 105 -250 155 -230
rect 105 -285 120 -250
rect 140 -285 155 -250
rect 105 -295 155 -285
rect 185 -195 235 -185
rect 185 -230 200 -195
rect 220 -230 235 -195
rect 185 -250 235 -230
rect 185 -285 200 -250
rect 220 -285 235 -250
rect 185 -295 235 -285
rect 250 -195 300 -185
rect 250 -230 265 -195
rect 285 -230 300 -195
rect 250 -250 300 -230
rect 250 -285 265 -250
rect 285 -285 300 -250
rect 250 -295 300 -285
rect 315 -195 360 -185
rect 315 -230 330 -195
rect 350 -230 360 -195
rect 315 -250 360 -230
rect 315 -285 330 -250
rect 350 -285 360 -250
rect 315 -295 360 -285
rect 435 -195 485 -185
rect 435 -230 450 -195
rect 470 -230 485 -195
rect 435 -250 485 -230
rect 435 -285 450 -250
rect 470 -285 485 -250
rect 435 -295 485 -285
rect 500 -195 545 -185
rect 500 -230 515 -195
rect 535 -230 545 -195
rect 500 -250 545 -230
rect 500 -285 515 -250
rect 535 -285 545 -250
rect 500 -295 545 -285
<< pdiff >>
rect -525 210 -475 220
rect -525 175 -510 210
rect -490 175 -475 210
rect -525 155 -475 175
rect -525 120 -510 155
rect -490 120 -475 155
rect -525 100 -475 120
rect -525 65 -510 100
rect -490 65 -475 100
rect -525 45 -475 65
rect -525 10 -510 45
rect -490 10 -475 45
rect -525 5 -475 10
rect -520 0 -475 5
rect -460 210 -410 220
rect -460 175 -445 210
rect -425 175 -410 210
rect -460 155 -410 175
rect -460 120 -445 155
rect -425 120 -410 155
rect -460 100 -410 120
rect -460 65 -445 100
rect -425 65 -410 100
rect -460 45 -410 65
rect -460 10 -445 45
rect -425 10 -410 45
rect -460 0 -410 10
rect -395 210 -350 220
rect -395 175 -380 210
rect -360 175 -350 210
rect -395 155 -350 175
rect -395 120 -380 155
rect -360 120 -350 155
rect -395 100 -350 120
rect -395 65 -380 100
rect -360 65 -350 100
rect -395 45 -350 65
rect -395 10 -380 45
rect -360 10 -350 45
rect -395 0 -350 10
rect -205 210 -160 220
rect -205 175 -195 210
rect -175 175 -160 210
rect -205 155 -160 175
rect -205 120 -195 155
rect -175 120 -160 155
rect -205 100 -160 120
rect -205 65 -195 100
rect -175 65 -160 100
rect -205 45 -160 65
rect -205 10 -195 45
rect -175 10 -160 45
rect -205 0 -160 10
rect -145 210 -95 220
rect -145 175 -130 210
rect -110 175 -95 210
rect -145 155 -95 175
rect -145 120 -130 155
rect -110 120 -95 155
rect -145 100 -95 120
rect -145 65 -130 100
rect -110 65 -95 100
rect -145 45 -95 65
rect -145 10 -130 45
rect -110 10 -95 45
rect -145 0 -95 10
rect -20 210 25 220
rect -20 175 -10 210
rect 10 175 25 210
rect -20 155 25 175
rect -20 120 -10 155
rect 10 120 25 155
rect -20 100 25 120
rect -20 65 -10 100
rect 10 65 25 100
rect -20 45 25 65
rect -20 10 -10 45
rect 10 10 25 45
rect -20 0 25 10
rect 40 210 90 220
rect 40 175 55 210
rect 75 175 90 210
rect 40 155 90 175
rect 40 120 55 155
rect 75 120 90 155
rect 40 100 90 120
rect 40 65 55 100
rect 75 65 90 100
rect 40 45 90 65
rect 40 10 55 45
rect 75 10 90 45
rect 40 0 90 10
rect 105 210 155 220
rect 105 175 120 210
rect 140 175 155 210
rect 105 155 155 175
rect 105 120 120 155
rect 140 120 155 155
rect 105 100 155 120
rect 105 65 120 100
rect 140 65 155 100
rect 105 45 155 65
rect 105 10 120 45
rect 140 10 155 45
rect 105 0 155 10
rect 185 210 235 220
rect 185 175 200 210
rect 220 175 235 210
rect 185 155 235 175
rect 185 120 200 155
rect 220 120 235 155
rect 185 100 235 120
rect 185 65 200 100
rect 220 65 235 100
rect 185 45 235 65
rect 185 10 200 45
rect 220 10 235 45
rect 185 0 235 10
rect 250 210 300 220
rect 250 175 265 210
rect 285 175 300 210
rect 250 155 300 175
rect 250 120 265 155
rect 285 120 300 155
rect 250 100 300 120
rect 250 65 265 100
rect 285 65 300 100
rect 250 45 300 65
rect 250 10 265 45
rect 285 10 300 45
rect 250 0 300 10
rect 315 210 360 220
rect 315 175 330 210
rect 350 175 360 210
rect 315 155 360 175
rect 315 120 330 155
rect 350 120 360 155
rect 315 100 360 120
rect 315 65 330 100
rect 350 65 360 100
rect 315 45 360 65
rect 315 10 330 45
rect 350 10 360 45
rect 315 0 360 10
rect 435 210 485 220
rect 435 175 450 210
rect 470 175 485 210
rect 435 155 485 175
rect 435 120 450 155
rect 470 120 485 155
rect 435 100 485 120
rect 435 65 450 100
rect 470 65 485 100
rect 435 45 485 65
rect 435 10 450 45
rect 470 10 485 45
rect 435 0 485 10
rect 500 210 545 220
rect 500 175 515 210
rect 535 175 545 210
rect 500 155 545 175
rect 500 120 515 155
rect 535 120 545 155
rect 500 100 545 120
rect 500 65 515 100
rect 535 65 545 100
rect 500 45 545 65
rect 500 10 515 45
rect 535 10 545 45
rect 500 0 545 10
<< ndiffc >>
rect -215 -230 -195 -195
rect -510 -285 -490 -250
rect -445 -285 -425 -250
rect -380 -285 -360 -250
rect -215 -285 -195 -250
rect -150 -230 -130 -195
rect -150 -285 -130 -250
rect -10 -230 10 -195
rect -10 -285 10 -250
rect 55 -230 75 -195
rect 55 -285 75 -250
rect 120 -230 140 -195
rect 120 -285 140 -250
rect 200 -230 220 -195
rect 200 -285 220 -250
rect 265 -230 285 -195
rect 265 -285 285 -250
rect 330 -230 350 -195
rect 330 -285 350 -250
rect 450 -230 470 -195
rect 450 -285 470 -250
rect 515 -230 535 -195
rect 515 -285 535 -250
<< pdiffc >>
rect -510 175 -490 210
rect -510 120 -490 155
rect -510 65 -490 100
rect -510 10 -490 45
rect -445 175 -425 210
rect -445 120 -425 155
rect -445 65 -425 100
rect -445 10 -425 45
rect -380 175 -360 210
rect -380 120 -360 155
rect -380 65 -360 100
rect -380 10 -360 45
rect -195 175 -175 210
rect -195 120 -175 155
rect -195 65 -175 100
rect -195 10 -175 45
rect -130 175 -110 210
rect -130 120 -110 155
rect -130 65 -110 100
rect -130 10 -110 45
rect -10 175 10 210
rect -10 120 10 155
rect -10 65 10 100
rect -10 10 10 45
rect 55 175 75 210
rect 55 120 75 155
rect 55 65 75 100
rect 55 10 75 45
rect 120 175 140 210
rect 120 120 140 155
rect 120 65 140 100
rect 120 10 140 45
rect 200 175 220 210
rect 200 120 220 155
rect 200 65 220 100
rect 200 10 220 45
rect 265 175 285 210
rect 265 120 285 155
rect 265 65 285 100
rect 265 10 285 45
rect 330 175 350 210
rect 330 120 350 155
rect 330 65 350 100
rect 330 10 350 45
rect 450 175 470 210
rect 450 120 470 155
rect 450 65 470 100
rect 450 10 470 45
rect 515 175 535 210
rect 515 120 535 155
rect 515 65 535 100
rect 515 10 535 45
<< psubdiff >>
rect -270 -195 -225 -185
rect -270 -230 -255 -195
rect -235 -230 -225 -195
rect -350 -250 -305 -240
rect -350 -285 -340 -250
rect -320 -285 -305 -250
rect -350 -295 -305 -285
rect -270 -250 -225 -230
rect -270 -285 -255 -250
rect -235 -285 -225 -250
rect -270 -295 -225 -285
rect -85 -195 -25 -185
rect -85 -230 -70 -195
rect -50 -230 -25 -195
rect -85 -250 -25 -230
rect -85 -285 -70 -250
rect -50 -285 -25 -250
rect -85 -295 -25 -285
rect 360 -195 405 -185
rect 360 -230 370 -195
rect 390 -230 405 -195
rect 360 -250 405 -230
rect 360 -285 370 -250
rect 390 -285 405 -250
rect 360 -295 405 -285
rect 545 -195 590 -185
rect 545 -230 555 -195
rect 575 -230 590 -195
rect 545 -250 590 -230
rect 545 -285 555 -250
rect 575 -285 590 -250
rect 545 -295 590 -285
<< nsubdiff >>
rect -350 210 -305 220
rect -350 175 -340 210
rect -320 175 -305 210
rect -350 155 -305 175
rect -350 120 -340 155
rect -320 120 -305 155
rect -350 100 -305 120
rect -350 65 -340 100
rect -320 65 -305 100
rect -350 45 -305 65
rect -350 10 -340 45
rect -320 10 -305 45
rect -350 0 -305 10
rect -250 210 -205 220
rect -250 175 -235 210
rect -215 175 -205 210
rect -250 155 -205 175
rect -250 120 -235 155
rect -215 120 -205 155
rect -250 100 -205 120
rect -250 65 -235 100
rect -215 65 -205 100
rect -250 45 -205 65
rect -250 10 -235 45
rect -215 10 -205 45
rect -250 0 -205 10
rect -65 210 -20 220
rect -65 175 -50 210
rect -30 175 -20 210
rect -65 155 -20 175
rect -65 120 -50 155
rect -30 120 -20 155
rect -65 100 -20 120
rect -65 65 -50 100
rect -30 65 -20 100
rect -65 45 -20 65
rect -65 10 -50 45
rect -30 10 -20 45
rect -65 0 -20 10
rect 360 210 405 220
rect 360 175 370 210
rect 390 175 405 210
rect 360 155 405 175
rect 360 120 370 155
rect 390 120 405 155
rect 360 100 405 120
rect 360 65 370 100
rect 390 65 405 100
rect 360 45 405 65
rect 360 10 370 45
rect 390 10 405 45
rect 360 0 405 10
rect 545 210 590 220
rect 545 175 555 210
rect 575 175 590 210
rect 545 155 590 175
rect 545 120 555 155
rect 575 120 590 155
rect 545 100 590 120
rect 545 65 555 100
rect 575 65 590 100
rect 545 45 590 65
rect 545 10 555 45
rect 575 10 590 45
rect 545 0 590 10
<< psubdiffcont >>
rect -255 -230 -235 -195
rect -340 -285 -320 -250
rect -255 -285 -235 -250
rect -70 -230 -50 -195
rect -70 -285 -50 -250
rect 370 -230 390 -195
rect 370 -285 390 -250
rect 555 -230 575 -195
rect 555 -285 575 -250
<< nsubdiffcont >>
rect -340 175 -320 210
rect -340 120 -320 155
rect -340 65 -320 100
rect -340 10 -320 45
rect -235 175 -215 210
rect -235 120 -215 155
rect -235 65 -215 100
rect -235 10 -215 45
rect -50 175 -30 210
rect -50 120 -30 155
rect -50 65 -30 100
rect -50 10 -30 45
rect 370 175 390 210
rect 370 120 390 155
rect 370 65 390 100
rect 370 10 390 45
rect 555 175 575 210
rect 555 120 575 155
rect 555 65 575 100
rect 555 10 575 45
<< poly >>
rect -160 260 250 275
rect -475 220 -460 235
rect -410 220 -395 235
rect -160 220 -145 260
rect 25 220 40 235
rect 90 220 105 235
rect 235 220 250 260
rect 300 220 315 235
rect 485 220 500 235
rect -475 -80 -460 0
rect -410 -20 -395 0
rect -410 -30 -370 -20
rect -410 -50 -400 -30
rect -380 -50 -370 -30
rect -410 -60 -370 -50
rect -475 -90 -435 -80
rect -475 -110 -465 -90
rect -445 -110 -435 -90
rect -475 -120 -435 -110
rect -475 -240 -460 -120
rect -410 -240 -395 -60
rect -160 -105 -145 0
rect -180 -120 -145 -105
rect -180 -185 -165 -120
rect 25 -185 40 0
rect 90 -20 105 0
rect 65 -30 105 -20
rect 65 -50 75 -30
rect 95 -50 105 -30
rect 65 -60 105 -50
rect 90 -185 105 -60
rect 235 -185 250 0
rect 300 -20 315 0
rect 300 -30 340 -20
rect 300 -50 310 -30
rect 330 -50 340 -30
rect 300 -60 340 -50
rect 300 -185 315 -60
rect 485 -185 500 0
rect -475 -310 -460 -295
rect -410 -310 -395 -295
rect -180 -310 -165 -295
rect 25 -335 40 -295
rect 90 -310 105 -295
rect 235 -310 250 -295
rect 300 -310 315 -295
rect 485 -335 500 -295
rect 25 -350 500 -335
<< polycont >>
rect -400 -50 -380 -30
rect -465 -110 -445 -90
rect 75 -50 95 -30
rect 310 -50 330 -30
<< locali >>
rect -390 275 -350 285
rect -390 255 -380 275
rect -360 255 -350 275
rect -390 220 -350 255
rect -205 275 -165 285
rect -205 255 -195 275
rect -175 255 -165 275
rect -205 220 -165 255
rect -20 275 20 285
rect -20 255 -10 275
rect 10 255 20 275
rect -20 220 20 255
rect 320 275 360 285
rect 320 255 330 275
rect 350 255 360 275
rect 320 220 360 255
rect 505 275 545 285
rect 505 255 515 275
rect 535 255 545 275
rect 505 220 545 255
rect -520 210 -480 220
rect -520 175 -510 210
rect -490 175 -480 210
rect -520 155 -480 175
rect -520 120 -510 155
rect -490 120 -480 155
rect -520 100 -480 120
rect -520 65 -510 100
rect -490 65 -480 100
rect -520 45 -480 65
rect -520 10 -510 45
rect -490 10 -480 45
rect -520 0 -480 10
rect -455 210 -415 220
rect -455 175 -445 210
rect -425 175 -415 210
rect -455 155 -415 175
rect -455 120 -445 155
rect -425 120 -415 155
rect -455 100 -415 120
rect -455 65 -445 100
rect -425 65 -415 100
rect -455 45 -415 65
rect -455 10 -445 45
rect -425 10 -415 45
rect -455 0 -415 10
rect -390 210 -310 220
rect -390 175 -380 210
rect -360 175 -340 210
rect -320 175 -310 210
rect -390 155 -310 175
rect -390 120 -380 155
rect -360 120 -340 155
rect -320 120 -310 155
rect -390 100 -310 120
rect -390 65 -380 100
rect -360 65 -340 100
rect -320 65 -310 100
rect -390 45 -310 65
rect -390 10 -380 45
rect -360 10 -340 45
rect -320 10 -310 45
rect -390 0 -310 10
rect -245 210 -165 220
rect -245 175 -235 210
rect -215 175 -195 210
rect -175 175 -165 210
rect -245 155 -165 175
rect -245 120 -235 155
rect -215 120 -195 155
rect -175 120 -165 155
rect -245 100 -165 120
rect -245 65 -235 100
rect -215 65 -195 100
rect -175 65 -165 100
rect -245 45 -165 65
rect -245 10 -235 45
rect -215 10 -195 45
rect -175 10 -165 45
rect -245 0 -165 10
rect -140 210 -100 220
rect -140 175 -130 210
rect -110 175 -100 210
rect -140 155 -100 175
rect -140 120 -130 155
rect -110 120 -100 155
rect -140 100 -100 120
rect -140 65 -130 100
rect -110 65 -100 100
rect -140 45 -100 65
rect -140 10 -130 45
rect -110 10 -100 45
rect -520 -140 -495 0
rect -140 -20 -100 10
rect -60 210 20 220
rect -60 175 -50 210
rect -30 175 -10 210
rect 10 175 20 210
rect -60 155 20 175
rect -60 120 -50 155
rect -30 120 -10 155
rect 10 120 20 155
rect -60 100 20 120
rect -60 65 -50 100
rect -30 65 -10 100
rect 10 65 20 100
rect -60 45 20 65
rect -60 10 -50 45
rect -30 10 -10 45
rect 10 10 20 45
rect -60 0 20 10
rect 45 210 85 220
rect 45 175 55 210
rect 75 175 85 210
rect 45 155 85 175
rect 45 120 55 155
rect 75 120 85 155
rect 45 100 85 120
rect 45 65 55 100
rect 75 65 85 100
rect 45 45 85 65
rect 45 10 55 45
rect 75 10 85 45
rect 45 0 85 10
rect 110 210 150 220
rect 110 175 120 210
rect 140 175 150 210
rect 110 155 150 175
rect 110 120 120 155
rect 140 120 150 155
rect 110 100 150 120
rect 110 65 120 100
rect 140 65 150 100
rect 110 45 150 65
rect 110 10 120 45
rect 140 10 150 45
rect 110 0 150 10
rect -410 -30 105 -20
rect -410 -50 -400 -30
rect -380 -50 75 -30
rect 95 -50 105 -30
rect -410 -60 105 -50
rect -475 -90 -325 -80
rect -475 -110 -465 -90
rect -445 -110 -355 -90
rect -335 -110 -325 -90
rect -475 -120 -325 -110
rect -140 -125 -100 -60
rect 130 -80 150 0
rect 190 210 230 220
rect 190 175 200 210
rect 220 175 230 210
rect 190 155 230 175
rect 190 120 200 155
rect 220 120 230 155
rect 190 100 230 120
rect 190 65 200 100
rect 220 65 230 100
rect 190 45 230 65
rect 190 10 200 45
rect 220 10 230 45
rect 190 0 230 10
rect 255 210 295 220
rect 255 175 265 210
rect 285 175 295 210
rect 255 155 295 175
rect 255 120 265 155
rect 285 120 295 155
rect 255 100 295 120
rect 255 65 265 100
rect 285 65 295 100
rect 255 45 295 65
rect 255 10 265 45
rect 285 10 295 45
rect 255 0 295 10
rect 320 210 400 220
rect 320 175 330 210
rect 350 175 370 210
rect 390 175 400 210
rect 320 155 400 175
rect 320 120 330 155
rect 350 120 370 155
rect 390 120 400 155
rect 320 100 400 120
rect 320 65 330 100
rect 350 65 370 100
rect 390 65 400 100
rect 320 45 400 65
rect 320 10 330 45
rect 350 10 370 45
rect 390 10 400 45
rect 320 0 400 10
rect 440 210 480 220
rect 440 175 450 210
rect 470 175 480 210
rect 440 155 480 175
rect 440 120 450 155
rect 470 120 480 155
rect 440 100 480 120
rect 440 65 450 100
rect 470 65 480 100
rect 440 45 480 65
rect 440 10 450 45
rect 470 10 480 45
rect 190 -80 210 0
rect 440 -20 480 10
rect 505 210 585 220
rect 505 175 515 210
rect 535 175 555 210
rect 575 175 585 210
rect 505 155 585 175
rect 505 120 515 155
rect 535 120 555 155
rect 575 120 585 155
rect 505 100 585 120
rect 505 65 515 100
rect 535 65 555 100
rect 575 65 585 100
rect 505 45 585 65
rect 505 10 515 45
rect 535 10 555 45
rect 575 10 585 45
rect 505 0 585 10
rect 300 -30 480 -20
rect 300 -50 310 -30
rect 330 -50 480 -30
rect 300 -60 480 -50
rect -520 -180 -415 -140
rect -520 -250 -480 -240
rect -520 -285 -510 -250
rect -490 -285 -480 -250
rect -520 -325 -480 -285
rect -455 -250 -415 -180
rect -160 -160 -100 -125
rect 45 -120 210 -80
rect 355 -90 395 -60
rect 355 -110 365 -90
rect 385 -110 395 -90
rect 355 -120 395 -110
rect -20 -150 20 -140
rect -265 -195 -185 -185
rect -265 -230 -255 -195
rect -235 -230 -215 -195
rect -195 -230 -185 -195
rect -455 -285 -445 -250
rect -425 -285 -415 -250
rect -455 -295 -415 -285
rect -390 -250 -310 -240
rect -390 -285 -380 -250
rect -360 -285 -340 -250
rect -320 -285 -310 -250
rect -390 -295 -310 -285
rect -265 -250 -185 -230
rect -265 -285 -255 -250
rect -235 -285 -215 -250
rect -195 -285 -185 -250
rect -265 -295 -185 -285
rect -160 -195 -120 -160
rect -20 -170 -10 -150
rect 10 -170 20 -150
rect -160 -230 -150 -195
rect -130 -230 -120 -195
rect -160 -250 -120 -230
rect -160 -285 -150 -250
rect -130 -285 -120 -250
rect -160 -295 -120 -285
rect -80 -195 -40 -185
rect -80 -230 -70 -195
rect -50 -230 -40 -195
rect -80 -250 -40 -230
rect -80 -285 -70 -250
rect -50 -285 -40 -250
rect -520 -345 -510 -325
rect -490 -345 -480 -325
rect -520 -355 -480 -345
rect -390 -325 -350 -295
rect -390 -345 -380 -325
rect -360 -345 -350 -325
rect -390 -355 -350 -345
rect -225 -325 -185 -295
rect -225 -345 -215 -325
rect -195 -345 -185 -325
rect -225 -355 -185 -345
rect -80 -325 -40 -285
rect -20 -195 20 -170
rect -20 -230 -10 -195
rect 10 -230 20 -195
rect -20 -250 20 -230
rect -20 -285 -10 -250
rect 10 -285 20 -250
rect -20 -295 20 -285
rect 45 -195 85 -120
rect 45 -230 55 -195
rect 75 -230 85 -195
rect 45 -250 85 -230
rect 45 -285 55 -250
rect 75 -285 85 -250
rect 45 -295 85 -285
rect 110 -150 150 -140
rect 110 -170 120 -150
rect 140 -170 150 -150
rect 110 -195 150 -170
rect 255 -150 295 -140
rect 255 -170 265 -150
rect 285 -170 295 -150
rect 110 -230 120 -195
rect 140 -230 150 -195
rect 110 -250 150 -230
rect 110 -285 120 -250
rect 140 -285 150 -250
rect 110 -295 150 -285
rect 190 -195 230 -185
rect 190 -230 200 -195
rect 220 -230 230 -195
rect 190 -250 230 -230
rect 190 -285 200 -250
rect 220 -285 230 -250
rect -80 -345 -70 -325
rect -50 -345 -40 -325
rect -80 -355 -40 -345
rect 190 -325 230 -285
rect 255 -195 295 -170
rect 255 -230 265 -195
rect 285 -230 295 -195
rect 255 -250 295 -230
rect 255 -285 265 -250
rect 285 -285 295 -250
rect 255 -295 295 -285
rect 320 -195 400 -185
rect 320 -230 330 -195
rect 350 -230 370 -195
rect 390 -230 400 -195
rect 320 -250 400 -230
rect 320 -285 330 -250
rect 350 -285 370 -250
rect 390 -285 400 -250
rect 320 -295 400 -285
rect 440 -195 480 -60
rect 440 -230 450 -195
rect 470 -230 480 -195
rect 440 -250 480 -230
rect 440 -285 450 -250
rect 470 -285 480 -250
rect 440 -295 480 -285
rect 505 -195 585 -185
rect 505 -230 515 -195
rect 535 -230 555 -195
rect 575 -230 585 -195
rect 505 -250 585 -230
rect 505 -285 515 -250
rect 535 -285 555 -250
rect 575 -285 585 -250
rect 505 -295 585 -285
rect 190 -345 200 -325
rect 220 -345 230 -325
rect 190 -355 230 -345
rect 320 -325 360 -295
rect 320 -345 330 -325
rect 350 -345 360 -325
rect 320 -355 360 -345
rect 505 -325 545 -295
rect 505 -345 515 -325
rect 535 -345 545 -325
rect 505 -355 545 -345
<< viali >>
rect -380 255 -360 275
rect -195 255 -175 275
rect -10 255 10 275
rect 330 255 350 275
rect 515 255 535 275
rect -355 -110 -335 -90
rect 365 -110 385 -90
rect -10 -170 10 -150
rect -510 -345 -490 -325
rect -380 -345 -360 -325
rect -215 -345 -195 -325
rect 120 -170 140 -150
rect 265 -170 285 -150
rect -70 -345 -50 -325
rect 200 -345 220 -325
rect 330 -345 350 -325
rect 515 -345 535 -325
<< metal1 >>
rect -545 275 610 285
rect -545 255 -380 275
rect -360 255 -195 275
rect -175 255 -10 275
rect 10 255 330 275
rect 350 255 515 275
rect 535 255 610 275
rect -545 245 610 255
rect -365 -90 395 -80
rect -365 -110 -355 -90
rect -335 -110 365 -90
rect 385 -110 395 -90
rect -365 -120 395 -110
rect -20 -150 295 -140
rect -20 -170 -10 -150
rect 10 -170 120 -150
rect 140 -170 265 -150
rect 285 -170 295 -150
rect -20 -175 295 -170
rect -545 -325 610 -315
rect -545 -345 -510 -325
rect -490 -345 -380 -325
rect -360 -345 -215 -325
rect -195 -345 -70 -325
rect -50 -345 200 -325
rect 220 -345 330 -325
rect 350 -345 515 -325
rect 535 -345 610 -325
rect -545 -355 610 -345
<< labels >>
flabel metal1 410 260 420 270 0 FreeSans 160 0 164 104 VDD
port 11 nsew
flabel metal1 -145 -345 -135 -335 0 FreeSans 160 0 -58 -120 GND
port 13 nsew
flabel poly 490 -120 500 -105 0 FreeSans 160 0 172 -30 A
port 7 nsew
flabel poly -160 -120 -150 -105 0 FreeSans 160 0 -32 -30 B
port 5 nsew
flabel locali 125 -105 130 -100 0 FreeSans 160 0 50 -42 SUM_OUT
port 14 nsew
flabel locali -490 -170 -485 -165 0 FreeSans 160 0 -196 -68 CARRY_OUT
port 15 nsew
<< end >>
