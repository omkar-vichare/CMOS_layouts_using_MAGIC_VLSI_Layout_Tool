magic
tech sky130A
timestamp 1734865608
<< nwell >>
rect -100 25 170 175
<< nmos >>
rect 20 -155 35 -45
rect 85 -155 100 -45
<< pmos >>
rect 20 45 35 155
rect 85 45 100 155
<< ndiff >>
rect -30 -55 20 -45
rect -30 -90 -15 -55
rect 5 -90 20 -55
rect -30 -110 20 -90
rect -30 -145 -15 -110
rect 5 -145 20 -110
rect -30 -155 20 -145
rect 35 -55 85 -45
rect 35 -90 50 -55
rect 70 -90 85 -55
rect 35 -110 85 -90
rect 35 -145 50 -110
rect 70 -145 85 -110
rect 35 -155 85 -145
rect 100 -55 150 -45
rect 100 -90 115 -55
rect 135 -90 150 -55
rect 100 -110 150 -90
rect 100 -145 115 -110
rect 135 -145 150 -110
rect 100 -155 150 -145
<< pdiff >>
rect -30 145 20 155
rect -30 110 -15 145
rect 5 110 20 145
rect -30 90 20 110
rect -30 55 -15 90
rect 5 55 20 90
rect -30 45 20 55
rect 35 145 85 155
rect 35 110 50 145
rect 70 110 85 145
rect 35 90 85 110
rect 35 55 50 90
rect 70 55 85 90
rect 35 45 85 55
rect 100 145 150 155
rect 100 110 115 145
rect 135 110 150 145
rect 100 90 150 110
rect 100 55 115 90
rect 135 55 150 90
rect 100 45 150 55
<< ndiffc >>
rect -15 -90 5 -55
rect -15 -145 5 -110
rect 50 -90 70 -55
rect 50 -145 70 -110
rect 115 -90 135 -55
rect 115 -145 135 -110
<< pdiffc >>
rect -15 110 5 145
rect -15 55 5 90
rect 50 110 70 145
rect 50 55 70 90
rect 115 110 135 145
rect 115 55 135 90
<< psubdiff >>
rect -80 -55 -30 -45
rect -80 -90 -65 -55
rect -40 -90 -30 -55
rect -80 -110 -30 -90
rect -80 -145 -65 -110
rect -40 -145 -30 -110
rect -80 -155 -30 -145
<< nsubdiff >>
rect -80 145 -30 155
rect -80 110 -65 145
rect -40 110 -30 145
rect -80 90 -30 110
rect -80 55 -65 90
rect -40 55 -30 90
rect -80 45 -30 55
<< psubdiffcont >>
rect -65 -90 -40 -55
rect -65 -145 -40 -110
<< nsubdiffcont >>
rect -65 110 -40 145
rect -65 55 -40 90
<< poly >>
rect 20 155 35 170
rect 85 155 100 170
rect 20 -45 35 45
rect 85 -45 100 45
rect 20 -170 35 -155
rect 85 -170 100 -155
<< locali >>
rect -25 205 15 210
rect -25 185 -15 205
rect 5 185 15 205
rect -25 155 15 185
rect 105 205 145 210
rect 105 185 115 205
rect 135 185 145 205
rect -75 145 15 155
rect -75 110 -65 145
rect -40 110 -15 145
rect 5 110 15 145
rect -75 90 15 110
rect -75 55 -65 90
rect -40 55 -15 90
rect 5 55 15 90
rect -75 45 15 55
rect 40 145 80 155
rect 40 110 50 145
rect 70 110 80 145
rect 40 90 80 110
rect 40 55 50 90
rect 70 55 80 90
rect 40 25 80 55
rect 105 145 145 185
rect 105 110 115 145
rect 135 110 145 145
rect 105 90 145 110
rect 105 55 115 90
rect 135 55 145 90
rect 105 45 145 55
rect 40 -15 145 25
rect -75 -55 15 -45
rect -75 -90 -65 -55
rect -40 -90 -15 -55
rect 5 -90 15 -55
rect -75 -110 15 -90
rect -75 -145 -65 -110
rect -40 -145 -15 -110
rect 5 -145 15 -110
rect -75 -155 15 -145
rect 40 -55 80 -45
rect 40 -90 50 -55
rect 70 -90 80 -55
rect 40 -110 80 -90
rect 40 -145 50 -110
rect 70 -145 80 -110
rect 40 -155 80 -145
rect 105 -55 145 -15
rect 105 -90 115 -55
rect 135 -90 145 -55
rect 105 -110 145 -90
rect 105 -145 115 -110
rect 135 -145 145 -110
rect 105 -155 145 -145
rect -25 -185 15 -155
rect -25 -205 -15 -185
rect 5 -205 15 -185
rect -25 -210 15 -205
<< viali >>
rect -15 185 5 205
rect 115 185 135 205
rect -15 -205 5 -185
<< metal1 >>
rect -100 205 170 210
rect -100 185 -15 205
rect 5 185 115 205
rect 135 185 170 205
rect -100 180 170 185
rect -105 -185 170 -180
rect -105 -205 -15 -185
rect 5 -205 170 -185
rect -105 -210 170 -205
<< labels >>
flabel poly 25 -30 30 -25 0 FreeSans 80 0 10 -12 A
port 2 nsew
flabel poly 90 -30 95 -25 0 FreeSans 80 0 36 -12 B
port 3 nsew
flabel locali 130 5 140 15 0 FreeSans 80 0 52 2 NAND_OUT
port 4 nsew
flabel metal1 50 190 60 200 0 FreeSans 80 0 20 76 VDD
port 5 nsew
flabel metal1 50 -200 60 -190 0 FreeSans 80 0 20 -8 GND
port 6 nsew
<< end >>
