*nand2gate_magic.cir

.include nand2_layout.spice

Xnand A B NAND_OUT VDD GND nand2_layout

.end
