magic
tech sky130A
timestamp 1734872444
<< nwell >>
rect -205 285 90 545
<< nmos >>
rect -75 0 -60 115
rect -5 0 10 115
<< pmos >>
rect -75 305 -60 525
rect -5 305 10 525
<< ndiff >>
rect -130 105 -75 115
rect -130 70 -120 105
rect -90 70 -75 105
rect -130 45 -75 70
rect -130 10 -115 45
rect -85 10 -75 45
rect -130 0 -75 10
rect -60 105 -5 115
rect -60 70 -45 105
rect -20 70 -5 105
rect -60 45 -5 70
rect -60 10 -45 45
rect -20 10 -5 45
rect -60 0 -5 10
rect 10 105 70 115
rect 10 70 25 105
rect 55 70 70 105
rect 10 45 70 70
rect 10 10 25 45
rect 55 10 70 45
rect 10 0 70 10
<< pdiff >>
rect -130 515 -75 525
rect -130 480 -115 515
rect -95 480 -75 515
rect -130 460 -75 480
rect -130 425 -115 460
rect -95 425 -75 460
rect -130 405 -75 425
rect -130 370 -115 405
rect -95 370 -75 405
rect -130 350 -75 370
rect -130 315 -115 350
rect -95 315 -75 350
rect -130 305 -75 315
rect -60 515 -5 525
rect -60 480 -45 515
rect -20 480 -5 515
rect -60 460 -5 480
rect -60 425 -45 460
rect -20 425 -5 460
rect -60 405 -5 425
rect -60 370 -45 405
rect -20 370 -5 405
rect -60 350 -5 370
rect -60 315 -45 350
rect -20 315 -5 350
rect -60 305 -5 315
rect 10 515 70 525
rect 10 480 30 515
rect 50 480 70 515
rect 10 460 70 480
rect 10 425 30 460
rect 50 425 70 460
rect 10 405 70 425
rect 10 370 30 405
rect 50 370 70 405
rect 10 350 70 370
rect 10 315 30 350
rect 50 315 70 350
rect 10 305 70 315
<< ndiffc >>
rect -120 70 -90 105
rect -115 10 -85 45
rect -45 70 -20 105
rect -45 10 -20 45
rect 25 70 55 105
rect 25 10 55 45
<< pdiffc >>
rect -115 480 -95 515
rect -115 425 -95 460
rect -115 370 -95 405
rect -115 315 -95 350
rect -45 480 -20 515
rect -45 425 -20 460
rect -45 370 -20 405
rect -45 315 -20 350
rect 30 480 50 515
rect 30 425 50 460
rect 30 370 50 405
rect 30 315 50 350
<< psubdiff >>
rect -185 105 -130 115
rect -185 70 -170 105
rect -140 70 -130 105
rect -185 45 -130 70
rect -185 10 -170 45
rect -140 10 -130 45
rect -185 0 -130 10
<< nsubdiff >>
rect -185 515 -130 525
rect -185 480 -170 515
rect -140 480 -130 515
rect -185 460 -130 480
rect -185 425 -170 460
rect -140 425 -130 460
rect -185 405 -130 425
rect -185 370 -170 405
rect -140 370 -130 405
rect -185 350 -130 370
rect -185 315 -170 350
rect -140 315 -130 350
rect -185 305 -130 315
<< psubdiffcont >>
rect -170 70 -140 105
rect -170 10 -140 45
<< nsubdiffcont >>
rect -170 480 -140 515
rect -170 425 -140 460
rect -170 370 -140 405
rect -170 315 -140 350
<< poly >>
rect -75 525 -60 540
rect -5 525 10 540
rect -75 115 -60 305
rect -5 115 10 305
rect -75 -15 -60 0
rect -5 -15 10 0
<< locali >>
rect -130 580 -80 585
rect -130 555 -120 580
rect -90 555 -80 580
rect -130 525 -80 555
rect -180 515 -80 525
rect -180 480 -170 515
rect -140 480 -115 515
rect -95 480 -80 515
rect -180 460 -80 480
rect -180 425 -170 460
rect -140 425 -115 460
rect -95 425 -80 460
rect -180 405 -80 425
rect -180 370 -170 405
rect -140 370 -115 405
rect -95 370 -80 405
rect -180 350 -80 370
rect -180 315 -170 350
rect -140 315 -115 350
rect -95 315 -80 350
rect -180 305 -80 315
rect -55 515 -10 525
rect -55 480 -45 515
rect -20 480 -10 515
rect -55 460 -10 480
rect -55 425 -45 460
rect -20 425 -10 460
rect -55 405 -10 425
rect -55 370 -45 405
rect -20 370 -10 405
rect -55 350 -10 370
rect -55 315 -45 350
rect -20 315 -10 350
rect -55 305 -10 315
rect 15 515 65 525
rect 15 480 30 515
rect 50 480 65 515
rect 15 460 65 480
rect 15 425 30 460
rect 50 425 65 460
rect 15 405 65 425
rect 15 370 30 405
rect 50 370 65 405
rect 15 350 65 370
rect 15 315 30 350
rect 50 315 65 350
rect 15 225 65 315
rect -55 185 65 225
rect -180 105 -80 115
rect -180 70 -170 105
rect -140 70 -120 105
rect -90 70 -80 105
rect -180 45 -80 70
rect -180 10 -170 45
rect -140 10 -115 45
rect -85 10 -80 45
rect -180 0 -80 10
rect -55 105 -10 185
rect -55 70 -45 105
rect -20 70 -10 105
rect -55 45 -10 70
rect -55 10 -45 45
rect -20 10 -10 45
rect -55 0 -10 10
rect 15 105 65 115
rect 15 70 25 105
rect 55 70 65 105
rect 15 45 65 70
rect 15 10 25 45
rect 55 10 65 45
rect -180 -35 -130 0
rect -180 -60 -170 -35
rect -140 -60 -130 -35
rect -180 -65 -130 -60
rect 15 -35 65 10
rect 15 -60 25 -35
rect 55 -60 65 -35
rect 15 -65 65 -60
<< viali >>
rect -120 555 -90 580
rect -170 -60 -140 -35
rect 25 -60 55 -35
<< metal1 >>
rect -205 580 90 585
rect -205 555 -120 580
rect -90 555 90 580
rect -205 550 90 555
rect -205 -35 90 -30
rect -205 -60 -170 -35
rect -140 -60 25 -35
rect 55 -60 90 -35
rect -205 -65 90 -60
<< labels >>
flabel metal1 -5 560 10 575 0 FreeSans 160 0 -2 224 VDD
port 2 nsew
flabel metal1 -55 -55 -40 -40 0 FreeSans 160 0 -22 -22 GND
port 4 nsew
flabel locali 30 200 45 215 0 FreeSans 160 0 12 80 NOR_OUT
port 6 nsew
flabel poly -75 160 -60 175 7 FreeSans 160 0 -30 64 A
port 8 w
flabel poly -5 160 10 175 3 FreeSans 160 0 -2 64 B
port 11 e
<< end >>
